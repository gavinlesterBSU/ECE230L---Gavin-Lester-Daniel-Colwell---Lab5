module circuit_a(
    input A,
    input B,
    input C,
    input D,
    output Y

    // Declare inputs
    // Declare Y output
);
    assign Y = (~A & D);
    // Enter logic equation here

endmodule
